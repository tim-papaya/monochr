
module pll_usb (
	reset_reset,
	clk_clk);	

	input		reset_reset;
	input		clk_clk;
endmodule
