-- pll_usb.vhd

-- Generated using ACDS version 14.1 186 at 2020.01.24.17:15:23

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity pll_usb is
	port (
		clk_clk     : in  std_logic := '0'; --     clk.clk
		clk_out_clk : out std_logic;        -- clk_out.clk
		reset_reset : in  std_logic := '0'  --   reset.reset
	);
end entity pll_usb;

architecture rtl of pll_usb is
	component pll_usb_altpll_0 is
		port (
			clk       : in  std_logic                     := 'X';             -- clk
			reset     : in  std_logic                     := 'X';             -- reset
			read      : in  std_logic                     := 'X';             -- read
			write     : in  std_logic                     := 'X';             -- write
			address   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata  : out std_logic_vector(31 downto 0);                    -- readdata
			writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c2        : out std_logic;                                        -- clk
			areset    : in  std_logic                     := 'X';             -- export
			c1        : out std_logic;                                        -- export
			c0        : out std_logic;                                        -- export
			locked    : out std_logic;                                        -- export
			phasedone : out std_logic                                         -- export
		);
	end component pll_usb_altpll_0;

begin

	altpll_0 : component pll_usb_altpll_0
		port map (
			clk       => clk_clk,     --       inclk_interface.clk
			reset     => reset_reset, -- inclk_interface_reset.reset
			read      => open,        --             pll_slave.read
			write     => open,        --                      .write
			address   => open,        --                      .address
			readdata  => open,        --                      .readdata
			writedata => open,        --                      .writedata
			c2        => clk_out_clk, --                    c2.clk
			areset    => open,        --        areset_conduit.export
			c1        => open,        --            c1_conduit.export
			c0        => open,        --            c0_conduit.export
			locked    => open,        --        locked_conduit.export
			phasedone => open         --     phasedone_conduit.export
		);

end architecture rtl; -- of pll_usb
